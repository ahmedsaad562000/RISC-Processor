LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY ArithmaticPart IS
    generic (n: integer := 16);
    PORT (
        sel  : IN  std_logic_vector(1 downto 0);
        a, b : IN  std_logic_vector(n-1 downto 0);
        s    : OUT std_logic_vector(n-1 downto 0);
        cout : OUT std_logic
    );
END entity ;

ARCHITECTURE partaimp OF ArithmaticPart IS
    component select_adder IS
        generic (n: integer := 16);
        PORT (
            a, b : IN  std_logic_vector(n-1 downto 0);
            cin  : IN  std_logic;
            s    : OUT std_logic_vector(n-1 downto 0);
            cout : OUT std_logic
           );
    END component;

    signal inpb : std_logic_vector(n-1 downto 0);
    signal cin :   std_logic;
BEGIN
    
inpb <= b WHEN sel = "00"
ELSE x"0001" WHEN sel = "01"
ELSE (not x"0001") WHEN sel = "10"
ELSE (not b);
 
cin <= '0' WHEN sel(1) = '0'
 ELSE '1';

  f0: select_adder generic map(16) port map(a, inpb, cin,s, cout);
 
END partaimp;



