LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_Decode_stage IS
END tb_Decode_stage;

ARCHITECTURE tb_Decode_stage_arch OF tb_Decode_stage IS
    COMPONENT Decode_stage IS
        PORT (
            RST : IN STD_LOGIC;
            CLK : IN STD_LOGIC;
            RSRC1_ADD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            RSRC2_ADD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            RDST_ADD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            PC_PLUS_ONE_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            OP_CODE : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            CAT_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
            IMM_OR_INPUT : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            Write_back_Enable : IN STD_LOGIC;
            Write_back_value : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            Write_back_ADD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            FLAGS : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            SET_CLEAR : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
            PC_PLUS_ONE_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            Write_back : OUT STD_LOGIC;
            MEM_SRC : OUT STD_LOGIC;
            SP_INC : OUT STD_LOGIC;
            SP_DEC : OUT STD_LOGIC;
            MEM_WRITE : OUT STD_LOGIC;
            Out_Signal : OUT STD_LOGIC;
            CALL_Signal : OUT STD_LOGIC;
            ALU_Operation : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
            CIN_Signal : OUT STD_LOGIC;
            MEM_TO_REG : OUT STD_LOGIC;
            RSRC1_Value : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            RSRC2_Value : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            ALU_SRC : OUT STD_LOGIC;
            RSRC1_ADD_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
            RSRC2_ADD_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
            RDST_ADD_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
            IMM_OR_IN_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
        );
    END COMPONENT;
    SIGNAL RST_test : STD_LOGIC;
    SIGNAL CLK_test : STD_LOGIC;
    SIGNAL RSRC1_ADD_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL RSRC2_ADD_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL RDST_ADD_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL PC_PLUS_ONE_IN_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL OP_CODE_test : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL CAT_IN_test : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL IMM_OR_INPUT_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Write_back_Enable_test : STD_LOGIC;
    SIGNAL Write_back_value_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Write_back_ADD_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL FLAGS_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL SET_CLEAR_test : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL PC_PLUS_ONE_OUT_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Write_back_test : STD_LOGIC;
    SIGNAL MEM_SRC_test : STD_LOGIC;
    SIGNAL SP_INC_test : STD_LOGIC;
    SIGNAL SP_DEC_test : STD_LOGIC;
    SIGNAL MEM_WRITE_test : STD_LOGIC;
    SIGNAL Out_Signal_test : STD_LOGIC;
    SIGNAL CALL_Signal_test : STD_LOGIC;
    SIGNAL ALU_Operation_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL CIN_Signal_test : STD_LOGIC;
    SIGNAL MEM_TO_REG_test : STD_LOGIC;
    SIGNAL RSRC1_Value_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL RSRC2_Value_test : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL ALU_SRC_test : STD_LOGIC;
    SIGNAL RSRC1_ADD_OUT_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL RSRC2_ADD_OUT_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL RDST_ADD_OUT_test : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL IMM_OR_IN_OUT_test : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
    DECODE_STAGE_BOX : Decode_stage PORT MAP(
        RST_test, CLK_test, RSRC1_ADD_test, RSRC2_ADD_test, RDST_ADD_test,
        PC_PLUS_ONE_IN_test, OP_CODE_test, CAT_IN_test, IMM_OR_INPUT_test, Write_back_Enable_test, Write_back_value_test,
        Write_back_ADD_test, FLAGS_test, SET_CLEAR_test, PC_PLUS_ONE_OUT_test, Write_back_test, MEM_SRC_test, SP_INC_test,
        SP_DEC_test, MEM_WRITE_test, Out_Signal_test, CALL_Signal_test, ALU_Operation_test, CIN_Signal_test, MEM_TO_REG_test,
        RSRC1_Value_test, RSRC2_Value_test, ALU_SRC_test, RSRC1_ADD_OUT_test, RSRC2_ADD_OUT_test, RDST_ADD_OUT_test, IMM_OR_IN_OUT_test);

    PROCESS
	begin
        CLK_test <= '0';
        WAIT FOR 5 ns;
        CLK_test <= '1';
        WAIT FOR 5 ns;
    END PROCESS;

    Process
	begin 
    RST_test <= '1';
    wait for 10 ns;
    ---------------------------------------------------------------
    -------------- Increment Instruction -------------------------
    RST_test <= '0';
    RSRC1_ADD_test <= "000";
    RSRC2_ADD_test <= "001";
    RDST_ADD_test <= "010";
    PC_PLUS_ONE_IN_test <= x"0001";
    OP_CODE_test <= "01001";
    CAT_IN_test <= "10";
    IMM_OR_INPUT_test <= x"0002";
    Write_back_Enable_test <= '0';
    Write_back_value_test <= x"0000";
    Write_back_ADD_test <= "111";
    FLAGS_test <= "000";
    wait for 10 ns;
    ------------- POP instruction --------------------------------
    RSRC1_ADD_test <= "010";
    RSRC2_ADD_test <= "011";
    RDST_ADD_test <= "010";
    PC_PLUS_ONE_IN_test <= x"0001";
    OP_CODE_test <= "10100";
    CAT_IN_test <= "01";
    IMM_OR_INPUT_test <= x"0002";
    Write_back_Enable_test <= '0';
    Write_back_value_test <= x"0000";
    Write_back_ADD_test <= "111";
    FLAGS_test <= "000";
    wait for 10 ns;
    wait;
    End Process;

END ARCHITECTURE;